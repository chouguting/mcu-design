library verilog;
use verilog.vl_types.all;
entity tb_pipeline_calculate is
end tb_pipeline_calculate;
