library verilog;
use verilog.vl_types.all;
entity testbench_alu_7bits is
end testbench_alu_7bits;
