library verilog;
use verilog.vl_types.all;
entity tb_timer_clock is
end tb_timer_clock;
