library verilog;
use verilog.vl_types.all;
entity tb_controlled_counter is
end tb_controlled_counter;
