library verilog;
use verilog.vl_types.all;
entity testbench_bcd_counter is
end testbench_bcd_counter;
