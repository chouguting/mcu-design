library verilog;
use verilog.vl_types.all;
entity middle_test is
end middle_test;
