library verilog;
use verilog.vl_types.all;
entity tb_CPU is
end tb_CPU;
