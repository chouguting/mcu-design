library verilog;
use verilog.vl_types.all;
entity tb_acc_counter_adder is
end tb_acc_counter_adder;
