library verilog;
use verilog.vl_types.all;
entity tb_traffic_light is
end tb_traffic_light;
