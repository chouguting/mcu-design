module Stack (
    stack_out,
    stack_in,
    push,
    pop,
    reset,
    clk
);

//--------
    output[10:0] stack_out;
    input[10:0] stack_in;
    input push,pop,reset,clk;

//-------
    reg[3:0] stack_ptr;
    reg[10:0] stack[15:0];
    wire[10:0] stack_out;
    wire[3:0] stk_index;

    assign stk_index = stack_ptr + 1;
    assign stack_out = stack[stack_ptr[3:0]];

    always @(posedge clk) begin
        if(reset) begin
            stack_ptr <= 4'b1111;
        end else if(push) begin
            stack[stk_index[3:0]] <= stack_in;
            stack_ptr <= stack_ptr + 1;
            
        end else if(pop) begin
            stack_ptr <= stack_ptr - 1;
        end
    
    end

endmodule
